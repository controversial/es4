package snake_types is
  type direction is (NORTH, EAST, SOUTH, WEST, NONE);
end package;
