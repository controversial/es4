-- needs a in filename to go first alphabetically so that this definition is available for
-- subsequent files
package snake_types is
  type direction is (NORTH, EAST, SOUTH, WEST, NONE);
end package;
